module vuantum

fn main() {
	println('hey there')
}